module CPU
(
    input clk_i, 
    input rst_i
);

// TODO: Implement your CPU here

// Do not change the name of these module instances.
// Instruction_Memory Instruction_Memory(
//     .addr_i     (), 
//     .instr_o    ()
// );

// PC PC(
//     .clk_i      (),
//     .rst_i      (),
//     .pc_i       (),
//     .pc_o       ()
// );

// Registers Registers(
//     .clk_i      (),
//     .rst_i      (),
//     .RS1addr_i  (),
//     .RS2addr_i  (),
//     .RDaddr_i   (), 
//     .RDdata_i   (),
//     .RegWrite_i (), 
//     .RS1data_o  (), 
//     .RS2data_o  () 
// );


endmodule
